// soc_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                               //                        clk.clk
		output wire        hps_0_h2f_reset_reset_n,               //            hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, //               hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //                           .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //                           .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //                           .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //                           .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //                           .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //                           .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //                           .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //                           .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //                           .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //                           .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //                           .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //                           .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //                           .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,     //                           .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,     //                           .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,     //                           .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,     //                           .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,     //                           .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,     //                           .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //                           .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //                           .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //                           .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //                           .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //                           .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //                           .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //                           .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //                           .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //                           .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //                           .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //                           .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //                           .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //                           .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //                           .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //                           .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //                           .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //                           .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //                           .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,    //                           .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,   //                           .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,   //                           .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,    //                           .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //                           .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //                           .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //                           .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //                           .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,     //                           .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,     //                           .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //                           .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //                           .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,  //                           .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,  //                           .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  //                           .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  //                           .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  //                           .hps_io_gpio_inst_GPIO61
		output wire [9:0]  leds_0_external_connection_export,     // leds_0_external_connection.export
		output wire [14:0] memory_mem_a,                          //                     memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                           .mem_ba
		output wire        memory_mem_ck,                         //                           .mem_ck
		output wire        memory_mem_ck_n,                       //                           .mem_ck_n
		output wire        memory_mem_cke,                        //                           .mem_cke
		output wire        memory_mem_cs_n,                       //                           .mem_cs_n
		output wire        memory_mem_ras_n,                      //                           .mem_ras_n
		output wire        memory_mem_cas_n,                      //                           .mem_cas_n
		output wire        memory_mem_we_n,                       //                           .mem_we_n
		output wire        memory_mem_reset_n,                    //                           .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //                           .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //                           .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //                           .mem_dqs_n
		output wire        memory_mem_odt,                        //                           .mem_odt
		output wire [3:0]  memory_mem_dm,                         //                           .mem_dm
		input  wire        memory_oct_rzqin,                      //                           .oct_rzqin
		output wire        pll_0_outclk2_clk,                     //              pll_0_outclk2.clk
		input  wire        reset_reset_n,                         //                      reset.reset_n
		output wire [12:0] sdram_controller_0_wire_addr,          //    sdram_controller_0_wire.addr
		output wire [1:0]  sdram_controller_0_wire_ba,            //                           .ba
		output wire        sdram_controller_0_wire_cas_n,         //                           .cas_n
		output wire        sdram_controller_0_wire_cke,           //                           .cke
		output wire        sdram_controller_0_wire_cs_n,          //                           .cs_n
		inout  wire [15:0] sdram_controller_0_wire_dq,            //                           .dq
		output wire [1:0]  sdram_controller_0_wire_dqm,           //                           .dqm
		output wire        sdram_controller_0_wire_ras_n,         //                           .ras_n
		output wire        sdram_controller_0_wire_we_n           //                           .we_n
	);

	wire          pll_0_outclk0_clk;                                                                // pll_0:outclk_0 -> [hps_0:f2h_axi_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, irq_mapper_002:clk, jtag_uart:clk, leds_0:clk, lua_cpu_0:clock_sink_clk, mm_interconnect_0:pll_0_outclk0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller:clk, rst_controller_001:clk, rst_controller_004:clk, sysid:clock, sysid_qsys_0:clock]
	wire          pll_0_outclk1_clk;                                                                // pll_0:outclk_1 -> [mm_interconnect_0:pll_0_outclk1_clk, rst_controller_003:clk, sdram_controller_0:clk]
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_dataa;                               // nios2_gen2_0:A_ci_multi_dataa -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_dataa
	wire          nios2_gen2_0_custom_instruction_master_multi_writerc;                             // nios2_gen2_0:A_ci_multi_writerc -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_result;                              // nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_result -> nios2_gen2_0:A_ci_multi_result
	wire          nios2_gen2_0_custom_instruction_master_clk;                                       // nios2_gen2_0:A_ci_multi_clock -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_clk
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_datab;                               // nios2_gen2_0:A_ci_multi_datab -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_datab
	wire          nios2_gen2_0_custom_instruction_master_start;                                     // nios2_gen2_0:A_ci_multi_start -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_start
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_b;                                   // nios2_gen2_0:A_ci_multi_b -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_b
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_c;                                   // nios2_gen2_0:A_ci_multi_c -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_c
	wire          nios2_gen2_0_custom_instruction_master_reset_req;                                 // nios2_gen2_0:A_ci_multi_reset_req -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire          nios2_gen2_0_custom_instruction_master_done;                                      // nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_done -> nios2_gen2_0:A_ci_multi_done
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_a;                                   // nios2_gen2_0:A_ci_multi_a -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_a
	wire          nios2_gen2_0_custom_instruction_master_clk_en;                                    // nios2_gen2_0:A_ci_multi_clk_en -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_clken
	wire          nios2_gen2_0_custom_instruction_master_reset;                                     // nios2_gen2_0:A_ci_multi_reset -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_reset
	wire          nios2_gen2_0_custom_instruction_master_multi_readrb;                              // nios2_gen2_0:A_ci_multi_readrb -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_readrb
	wire          nios2_gen2_0_custom_instruction_master_multi_readra;                              // nios2_gen2_0:A_ci_multi_readra -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_readra
	wire    [7:0] nios2_gen2_0_custom_instruction_master_multi_n;                                   // nios2_gen2_0:A_ci_multi_n -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_n
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_readra -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire    [4:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a;              // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_a -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_a
	wire    [4:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b;              // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_b -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_b
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk;            // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_clk -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire    [4:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c;              // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_c -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_c
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start;          // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_start -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_start
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req;      // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done;           // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_done
	wire    [7:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n;              // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_n -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_n
	wire   [31:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_result
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_clken -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire   [31:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab;          // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_datab -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire   [31:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa;          // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset;          // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_reset -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire          nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc;        // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a;               // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b;               // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c;               // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk;             // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start;           // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req;       // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done;            // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_done
	wire    [7:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n;               // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result;          // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_result
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab;           // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa;           // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset;           // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire          nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_readra;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_readra -> lua_cpu_0:nios_lua_exec_slave_readra
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_a;       // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_a -> lua_cpu_0:nios_lua_exec_slave_a
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_b;       // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_b -> lua_cpu_0:nios_lua_exec_slave_b
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_readrb;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_readrb -> lua_cpu_0:nios_lua_exec_slave_readrb
	wire    [4:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_c;       // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_c -> lua_cpu_0:nios_lua_exec_slave_c
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk;     // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> lua_cpu_0:nios_lua_exec_slave_clk
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start;   // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> lua_cpu_0:nios_lua_exec_slave_start
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done;    // lua_cpu_0:nios_lua_exec_slave_done -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire    [1:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_n;       // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_n -> lua_cpu_0:nios_lua_exec_slave_n
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result;  // lua_cpu_0:nios_lua_exec_slave_result -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_clken -> lua_cpu_0:nios_lua_exec_slave_clk_en
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab;   // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_datab -> lua_cpu_0:nios_lua_exec_slave_datab
	wire   [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa;   // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> lua_cpu_0:nios_lua_exec_slave_dataa
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset;   // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> lua_cpu_0:nios_lua_exec_slave_reset
	wire          nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_writerc; // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_writerc -> lua_cpu_0:nios_lua_exec_slave_writerc
	wire   [31:0] lua_cpu_0_avalon_master_readdata;                                                 // mm_interconnect_0:lua_cpu_0_avalon_master_readdata -> lua_cpu_0:avalon_master_readdata
	wire          lua_cpu_0_avalon_master_waitrequest;                                              // mm_interconnect_0:lua_cpu_0_avalon_master_waitrequest -> lua_cpu_0:avalon_master_waitrequest
	wire   [31:0] lua_cpu_0_avalon_master_address;                                                  // lua_cpu_0:avalon_master_address -> mm_interconnect_0:lua_cpu_0_avalon_master_address
	wire          lua_cpu_0_avalon_master_read;                                                     // lua_cpu_0:avalon_master_read -> mm_interconnect_0:lua_cpu_0_avalon_master_read
	wire   [31:0] lua_cpu_0_avalon_master_writedata;                                                // lua_cpu_0:avalon_master_writedata -> mm_interconnect_0:lua_cpu_0_avalon_master_writedata
	wire          lua_cpu_0_avalon_master_write;                                                    // lua_cpu_0:avalon_master_write -> mm_interconnect_0:lua_cpu_0_avalon_master_write
	wire   [31:0] nios2_gen2_0_data_master_readdata;                                                // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire          nios2_gen2_0_data_master_waitrequest;                                             // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire          nios2_gen2_0_data_master_debugaccess;                                             // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire   [30:0] nios2_gen2_0_data_master_address;                                                 // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire    [3:0] nios2_gen2_0_data_master_byteenable;                                              // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire          nios2_gen2_0_data_master_read;                                                    // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire          nios2_gen2_0_data_master_write;                                                   // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire   [31:0] nios2_gen2_0_data_master_writedata;                                               // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [31:0] nios2_gen2_0_instruction_master_readdata;                                         // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire          nios2_gen2_0_instruction_master_waitrequest;                                      // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire   [30:0] nios2_gen2_0_instruction_master_address;                                          // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire          nios2_gen2_0_instruction_master_read;                                             // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire          nios2_gen2_0_instruction_master_readdatavalid;                                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                                     // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                                       // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                                       // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                                      // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                         // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                                      // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                                       // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                         // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                                     // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                                      // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                                      // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                                      // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                                      // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                                       // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                                     // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                                     // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                                        // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                                      // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                                      // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                                      // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                                       // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                                     // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                                       // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                                     // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                                     // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                                      // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                                      // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                                       // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                                       // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                                       // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                                        // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                         // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                                      // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                                      // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                                     // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                                      // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                                  // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                                    // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                                    // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                                   // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                                    // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                                      // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                                  // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                                   // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                                   // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                                   // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                                   // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                                    // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                                  // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                                  // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                                     // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                                   // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                                   // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                                   // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                                  // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                                   // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                                   // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                                    // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                                     // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                                   // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                                  // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire          mm_interconnect_0_sdram_controller_0_s1_chipselect;                               // mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	wire   [15:0] mm_interconnect_0_sdram_controller_0_s1_readdata;                                 // sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	wire          mm_interconnect_0_sdram_controller_0_s1_waitrequest;                              // sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	wire   [24:0] mm_interconnect_0_sdram_controller_0_s1_address;                                  // mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	wire          mm_interconnect_0_sdram_controller_0_s1_read;                                     // mm_interconnect_0:sdram_controller_0_s1_read -> sdram_controller_0:az_rd_n
	wire    [1:0] mm_interconnect_0_sdram_controller_0_s1_byteenable;                               // mm_interconnect_0:sdram_controller_0_s1_byteenable -> sdram_controller_0:az_be_n
	wire          mm_interconnect_0_sdram_controller_0_s1_readdatavalid;                            // sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	wire          mm_interconnect_0_sdram_controller_0_s1_write;                                    // mm_interconnect_0:sdram_controller_0_s1_write -> sdram_controller_0:az_wr_n
	wire   [15:0] mm_interconnect_0_sdram_controller_0_s1_writedata;                                // mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                          // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                       // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                            // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                             // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire          mm_interconnect_0_leds_0_s1_chipselect;                                           // mm_interconnect_0:leds_0_s1_chipselect -> leds_0:chipselect
	wire   [31:0] mm_interconnect_0_leds_0_s1_readdata;                                             // leds_0:readdata -> mm_interconnect_0:leds_0_s1_readdata
	wire    [1:0] mm_interconnect_0_leds_0_s1_address;                                              // mm_interconnect_0:leds_0_s1_address -> leds_0:address
	wire          mm_interconnect_0_leds_0_s1_write;                                                // mm_interconnect_0:leds_0_s1_write -> leds_0:write_n
	wire   [31:0] mm_interconnect_0_leds_0_s1_writedata;                                            // mm_interconnect_0:leds_0_s1_writedata -> leds_0:writedata
	wire   [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                   // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_control_slave_address;                                    // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                 // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [63:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire    [7:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                 // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                                      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [63:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                                      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire   [31:0] hps_0_f2h_irq0_irq;                                                               // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                               // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire   [31:0] nios2_gen2_0_irq_irq;                                                             // irq_mapper_002:sender_irq -> nios2_gen2_0:irq
	wire          irq_mapper_receiver0_irq;                                                         // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq]
	wire          rst_controller_reset_out_reset;                                                   // rst_controller:reset_out -> [irq_mapper_002:reset, jtag_uart:rst_n, leds_0:reset_n, lua_cpu_0:reset_sink_reset, mm_interconnect_0:lua_cpu_0_reset_sink_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, sysid:reset_n, sysid_qsys_0:reset_n]
	wire          rst_controller_reset_out_reset_req;                                               // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire          nios2_gen2_0_debug_reset_request_reset;                                           // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                               // rst_controller_001:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire          rst_controller_001_reset_out_reset_req;                                           // rst_controller_001:reset_req -> onchip_memory2_0:reset_req
	wire          rst_controller_002_reset_out_reset;                                               // rst_controller_002:reset_out -> pll_0:rst
	wire          rst_controller_003_reset_out_reset;                                               // rst_controller_003:reset_out -> [mm_interconnect_0:sdram_controller_0_reset_reset_bridge_in_reset_reset, sdram_controller_0:reset_n]
	wire          rst_controller_004_reset_out_reset;                                               // rst_controller_004:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                          //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                         //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                         //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                       //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                        //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                       //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                      //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                      //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                       //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                    //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                         //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                        //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                      //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                        //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                         //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                      //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),    //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),   //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),   //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),    //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),  //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),  //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),  //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),               //         h2f_reset.reset_n
		.h2f_axi_clk              (pll_0_outclk0_clk),                     //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),             //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),           //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),            //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),           //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),          //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),           //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),          //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),           //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),          //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),          //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),              //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),            //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),            //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),            //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),           //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),           //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),              //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),            //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),           //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),           //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),             //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),           //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),            //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),           //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),          //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),           //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),          //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),           //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),          //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),          //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),              //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),            //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),            //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),            //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),           //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),           //                  .rready
		.f2h_axi_clk              (pll_0_outclk0_clk),                     //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                      //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                      //                  .awaddr
		.f2h_AWLEN                (),                                      //                  .awlen
		.f2h_AWSIZE               (),                                      //                  .awsize
		.f2h_AWBURST              (),                                      //                  .awburst
		.f2h_AWLOCK               (),                                      //                  .awlock
		.f2h_AWCACHE              (),                                      //                  .awcache
		.f2h_AWPROT               (),                                      //                  .awprot
		.f2h_AWVALID              (),                                      //                  .awvalid
		.f2h_AWREADY              (),                                      //                  .awready
		.f2h_AWUSER               (),                                      //                  .awuser
		.f2h_WID                  (),                                      //                  .wid
		.f2h_WDATA                (),                                      //                  .wdata
		.f2h_WSTRB                (),                                      //                  .wstrb
		.f2h_WLAST                (),                                      //                  .wlast
		.f2h_WVALID               (),                                      //                  .wvalid
		.f2h_WREADY               (),                                      //                  .wready
		.f2h_BID                  (),                                      //                  .bid
		.f2h_BRESP                (),                                      //                  .bresp
		.f2h_BVALID               (),                                      //                  .bvalid
		.f2h_BREADY               (),                                      //                  .bready
		.f2h_ARID                 (),                                      //                  .arid
		.f2h_ARADDR               (),                                      //                  .araddr
		.f2h_ARLEN                (),                                      //                  .arlen
		.f2h_ARSIZE               (),                                      //                  .arsize
		.f2h_ARBURST              (),                                      //                  .arburst
		.f2h_ARLOCK               (),                                      //                  .arlock
		.f2h_ARCACHE              (),                                      //                  .arcache
		.f2h_ARPROT               (),                                      //                  .arprot
		.f2h_ARVALID              (),                                      //                  .arvalid
		.f2h_ARREADY              (),                                      //                  .arready
		.f2h_ARUSER               (),                                      //                  .aruser
		.f2h_RID                  (),                                      //                  .rid
		.f2h_RDATA                (),                                      //                  .rdata
		.f2h_RRESP                (),                                      //                  .rresp
		.f2h_RLAST                (),                                      //                  .rlast
		.f2h_RVALID               (),                                      //                  .rvalid
		.f2h_RREADY               (),                                      //                  .rready
		.h2f_lw_axi_clk           (pll_0_outclk0_clk),                     //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),        //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),         //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),        //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),       //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),        //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),       //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),        //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),       //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),       //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),           //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),         //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),         //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),         //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),        //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),        //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),           //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),         //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),        //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),        //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),          //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),        //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),         //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),        //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),       //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),        //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),       //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),        //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),       //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),       //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),           //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),         //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),         //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),         //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),        //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),        //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                    //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                     //          f2h_irq1.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (pll_0_outclk0_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	soc_system_leds_0 leds_0 (
		.clk        (pll_0_outclk0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_leds_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_0_s1_readdata),   //                    .readdata
		.out_port   (leds_0_external_connection_export)       // external_connection.export
	);

	soc_system_lua_cpu_0 lua_cpu_0 (
		.nios_lua_exec_slave_dataa   (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),   // nios_lua_exec_slave.dataa
		.nios_lua_exec_slave_datab   (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),   //                    .datab
		.nios_lua_exec_slave_result  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result),  //                    .result
		.nios_lua_exec_slave_clk     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),     //                    .clk
		.nios_lua_exec_slave_clk_en  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),  //                    .clk_en
		.nios_lua_exec_slave_start   (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start),   //                    .start
		.nios_lua_exec_slave_done    (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done),    //                    .done
		.nios_lua_exec_slave_a       (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_a),       //                    .a
		.nios_lua_exec_slave_b       (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_b),       //                    .b
		.nios_lua_exec_slave_c       (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_c),       //                    .c
		.nios_lua_exec_slave_n       (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_n),       //                    .n
		.nios_lua_exec_slave_readra  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_readra),  //                    .readra
		.nios_lua_exec_slave_readrb  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_readrb),  //                    .readrb
		.nios_lua_exec_slave_reset   (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),   //                    .reset
		.nios_lua_exec_slave_writerc (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_writerc), //                    .writerc
		.avalon_master_address       (lua_cpu_0_avalon_master_address),                                                  //       avalon_master.address
		.avalon_master_readdata      (lua_cpu_0_avalon_master_readdata),                                                 //                    .readdata
		.avalon_master_writedata     (lua_cpu_0_avalon_master_writedata),                                                //                    .writedata
		.avalon_master_read          (lua_cpu_0_avalon_master_read),                                                     //                    .read
		.avalon_master_write         (lua_cpu_0_avalon_master_write),                                                    //                    .write
		.avalon_master_waitrequest   (lua_cpu_0_avalon_master_waitrequest),                                              //                    .waitrequest
		.clock_sink_clk              (pll_0_outclk0_clk),                                                                //          clock_sink.clk
		.reset_sink_reset            (rst_controller_reset_out_reset)                                                    //          reset_sink.reset
	);

	soc_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_0_outclk0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_gen2_0_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_gen2_0_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_gen2_0_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_gen2_0_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_gen2_0_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_gen2_0_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_gen2_0_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_gen2_0_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_gen2_0_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_gen2_0_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_gen2_0_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_gen2_0_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_gen2_0_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_gen2_0_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_gen2_0_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_gen2_0_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	soc_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_0_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_system_pll_0 pll_0 (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_002_reset_out_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),                  // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk),                  // outclk1.clk
		.outclk_2 (pll_0_outclk2_clk),                  // outclk2.clk
		.locked   ()                                    // (terminated)
	);

	soc_system_sdram_controller_0 sdram_controller_0 (
		.clk            (pll_0_outclk1_clk),                                     //   clk.clk
		.reset_n        (~rst_controller_003_reset_out_reset),                   // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_0_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_0_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_0_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_0_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_0_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_0_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_0_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_0_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_0_wire_we_n)                           //      .export
	);

	soc_system_sysid sysid (
		.clock    (pll_0_outclk0_clk),                              //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	soc_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_0_outclk0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_gen2_0_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                            //        ci_slave.result
		.ci_slave_multi_clk        (nios2_gen2_0_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_gen2_0_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_gen2_0_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_gen2_0_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_gen2_0_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_gen2_0_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_gen2_0_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_gen2_0_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_gen2_0_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_gen2_0_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_gen2_0_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_gen2_0_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_gen2_0_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_gen2_0_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_gen2_0_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_gen2_0_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                            //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_n                (8'b00000000),                                                                 //     (terminated)
		.ci_slave_readra           (1'b0),                                                                        //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                        //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                        //     (terminated)
		.ci_slave_a                (5'b00000),                                                                    //     (terminated)
		.ci_slave_b                (5'b00000),                                                                    //     (terminated)
		.ci_slave_c                (5'b00000),                                                                    //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                        //     (terminated)
		.comb_ci_master_dataa      (),                                                                            //     (terminated)
		.comb_ci_master_datab      (),                                                                            //     (terminated)
		.comb_ci_master_n          (),                                                                            //     (terminated)
		.comb_ci_master_readra     (),                                                                            //     (terminated)
		.comb_ci_master_readrb     (),                                                                            //     (terminated)
		.comb_ci_master_writerc    (),                                                                            //     (terminated)
		.comb_ci_master_a          (),                                                                            //     (terminated)
		.comb_ci_master_b          (),                                                                            //     (terminated)
		.comb_ci_master_c          (),                                                                            //     (terminated)
		.comb_ci_master_ipending   (),                                                                            //     (terminated)
		.comb_ci_master_estatus    ()                                                                             //     (terminated)
	);

	soc_system_nios2_gen2_0_custom_instruction_master_multi_xconnect nios2_gen2_0_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                            //           .ipending
		.ci_slave_estatus     (),                                                                            //           .estatus
		.ci_slave_clk         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_gen2_0_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),           //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab),           //          .datab
		.ci_slave_result     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result),          //          .result
		.ci_slave_n          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n),               //          .n
		.ci_slave_readra     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra),          //          .readra
		.ci_slave_readrb     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),          //          .readrb
		.ci_slave_writerc    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),         //          .writerc
		.ci_slave_a          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a),               //          .a
		.ci_slave_b          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b),               //          .b
		.ci_slave_c          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c),               //          .c
		.ci_slave_ipending   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),        //          .ipending
		.ci_slave_estatus    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),         //          .estatus
		.ci_slave_clk        (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk),             //          .clk
		.ci_slave_clken      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),          //          .clk_en
		.ci_slave_reset_req  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),       //          .reset_req
		.ci_slave_reset      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset),           //          .reset
		.ci_slave_start      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start),           //          .start
		.ci_slave_done       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done),            //          .done
		.ci_master_dataa     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),   // ci_master.dataa
		.ci_master_datab     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),   //          .datab
		.ci_master_result    (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result),  //          .result
		.ci_master_n         (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_n),       //          .n
		.ci_master_readra    (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_readra),  //          .readra
		.ci_master_readrb    (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_readrb),  //          .readrb
		.ci_master_writerc   (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_writerc), //          .writerc
		.ci_master_a         (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_a),       //          .a
		.ci_master_b         (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_b),       //          .b
		.ci_master_c         (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_c),       //          .c
		.ci_master_clk       (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),     //          .clk
		.ci_master_clken     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),  //          .clk_en
		.ci_master_reset     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),   //          .reset
		.ci_master_start     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start),   //          .start
		.ci_master_done      (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done),    //          .done
		.ci_master_ipending  (),                                                                                 // (terminated)
		.ci_master_estatus   (),                                                                                 // (terminated)
		.ci_master_reset_req ()                                                                                  // (terminated)
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                  //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                 //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                               //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                               //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                               //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                               //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                   //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                 //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                 //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                 //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                   //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                 //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                  //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                 //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                               //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                               //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                               //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                               //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                   //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                 //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                 //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                 //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                //                                                           .rready
		.hps_0_h2f_lw_axi_master_awid                                     (hps_0_h2f_lw_axi_master_awid),                               //                                    hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                   (hps_0_h2f_lw_axi_master_awaddr),                             //                                                           .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                    (hps_0_h2f_lw_axi_master_awlen),                              //                                                           .awlen
		.hps_0_h2f_lw_axi_master_awsize                                   (hps_0_h2f_lw_axi_master_awsize),                             //                                                           .awsize
		.hps_0_h2f_lw_axi_master_awburst                                  (hps_0_h2f_lw_axi_master_awburst),                            //                                                           .awburst
		.hps_0_h2f_lw_axi_master_awlock                                   (hps_0_h2f_lw_axi_master_awlock),                             //                                                           .awlock
		.hps_0_h2f_lw_axi_master_awcache                                  (hps_0_h2f_lw_axi_master_awcache),                            //                                                           .awcache
		.hps_0_h2f_lw_axi_master_awprot                                   (hps_0_h2f_lw_axi_master_awprot),                             //                                                           .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                  (hps_0_h2f_lw_axi_master_awvalid),                            //                                                           .awvalid
		.hps_0_h2f_lw_axi_master_awready                                  (hps_0_h2f_lw_axi_master_awready),                            //                                                           .awready
		.hps_0_h2f_lw_axi_master_wid                                      (hps_0_h2f_lw_axi_master_wid),                                //                                                           .wid
		.hps_0_h2f_lw_axi_master_wdata                                    (hps_0_h2f_lw_axi_master_wdata),                              //                                                           .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                    (hps_0_h2f_lw_axi_master_wstrb),                              //                                                           .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                    (hps_0_h2f_lw_axi_master_wlast),                              //                                                           .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                   (hps_0_h2f_lw_axi_master_wvalid),                             //                                                           .wvalid
		.hps_0_h2f_lw_axi_master_wready                                   (hps_0_h2f_lw_axi_master_wready),                             //                                                           .wready
		.hps_0_h2f_lw_axi_master_bid                                      (hps_0_h2f_lw_axi_master_bid),                                //                                                           .bid
		.hps_0_h2f_lw_axi_master_bresp                                    (hps_0_h2f_lw_axi_master_bresp),                              //                                                           .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                   (hps_0_h2f_lw_axi_master_bvalid),                             //                                                           .bvalid
		.hps_0_h2f_lw_axi_master_bready                                   (hps_0_h2f_lw_axi_master_bready),                             //                                                           .bready
		.hps_0_h2f_lw_axi_master_arid                                     (hps_0_h2f_lw_axi_master_arid),                               //                                                           .arid
		.hps_0_h2f_lw_axi_master_araddr                                   (hps_0_h2f_lw_axi_master_araddr),                             //                                                           .araddr
		.hps_0_h2f_lw_axi_master_arlen                                    (hps_0_h2f_lw_axi_master_arlen),                              //                                                           .arlen
		.hps_0_h2f_lw_axi_master_arsize                                   (hps_0_h2f_lw_axi_master_arsize),                             //                                                           .arsize
		.hps_0_h2f_lw_axi_master_arburst                                  (hps_0_h2f_lw_axi_master_arburst),                            //                                                           .arburst
		.hps_0_h2f_lw_axi_master_arlock                                   (hps_0_h2f_lw_axi_master_arlock),                             //                                                           .arlock
		.hps_0_h2f_lw_axi_master_arcache                                  (hps_0_h2f_lw_axi_master_arcache),                            //                                                           .arcache
		.hps_0_h2f_lw_axi_master_arprot                                   (hps_0_h2f_lw_axi_master_arprot),                             //                                                           .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                  (hps_0_h2f_lw_axi_master_arvalid),                            //                                                           .arvalid
		.hps_0_h2f_lw_axi_master_arready                                  (hps_0_h2f_lw_axi_master_arready),                            //                                                           .arready
		.hps_0_h2f_lw_axi_master_rid                                      (hps_0_h2f_lw_axi_master_rid),                                //                                                           .rid
		.hps_0_h2f_lw_axi_master_rdata                                    (hps_0_h2f_lw_axi_master_rdata),                              //                                                           .rdata
		.hps_0_h2f_lw_axi_master_rresp                                    (hps_0_h2f_lw_axi_master_rresp),                              //                                                           .rresp
		.hps_0_h2f_lw_axi_master_rlast                                    (hps_0_h2f_lw_axi_master_rlast),                              //                                                           .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                   (hps_0_h2f_lw_axi_master_rvalid),                             //                                                           .rvalid
		.hps_0_h2f_lw_axi_master_rready                                   (hps_0_h2f_lw_axi_master_rready),                             //                                                           .rready
		.pll_0_outclk0_clk                                                (pll_0_outclk0_clk),                                          //                                              pll_0_outclk0.clk
		.pll_0_outclk1_clk                                                (pll_0_outclk1_clk),                                          //                                              pll_0_outclk1.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                         // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.lua_cpu_0_reset_sink_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                             //                 lua_cpu_0_reset_sink_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),                         //              onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.sdram_controller_0_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                         //             sdram_controller_0_reset_reset_bridge_in_reset.reset
		.lua_cpu_0_avalon_master_address                                  (lua_cpu_0_avalon_master_address),                            //                                    lua_cpu_0_avalon_master.address
		.lua_cpu_0_avalon_master_waitrequest                              (lua_cpu_0_avalon_master_waitrequest),                        //                                                           .waitrequest
		.lua_cpu_0_avalon_master_read                                     (lua_cpu_0_avalon_master_read),                               //                                                           .read
		.lua_cpu_0_avalon_master_readdata                                 (lua_cpu_0_avalon_master_readdata),                           //                                                           .readdata
		.lua_cpu_0_avalon_master_write                                    (lua_cpu_0_avalon_master_write),                              //                                                           .write
		.lua_cpu_0_avalon_master_writedata                                (lua_cpu_0_avalon_master_writedata),                          //                                                           .writedata
		.nios2_gen2_0_data_master_address                                 (nios2_gen2_0_data_master_address),                           //                                   nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                             (nios2_gen2_0_data_master_waitrequest),                       //                                                           .waitrequest
		.nios2_gen2_0_data_master_byteenable                              (nios2_gen2_0_data_master_byteenable),                        //                                                           .byteenable
		.nios2_gen2_0_data_master_read                                    (nios2_gen2_0_data_master_read),                              //                                                           .read
		.nios2_gen2_0_data_master_readdata                                (nios2_gen2_0_data_master_readdata),                          //                                                           .readdata
		.nios2_gen2_0_data_master_write                                   (nios2_gen2_0_data_master_write),                             //                                                           .write
		.nios2_gen2_0_data_master_writedata                               (nios2_gen2_0_data_master_writedata),                         //                                                           .writedata
		.nios2_gen2_0_data_master_debugaccess                             (nios2_gen2_0_data_master_debugaccess),                       //                                                           .debugaccess
		.nios2_gen2_0_instruction_master_address                          (nios2_gen2_0_instruction_master_address),                    //                            nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                      (nios2_gen2_0_instruction_master_waitrequest),                //                                                           .waitrequest
		.nios2_gen2_0_instruction_master_read                             (nios2_gen2_0_instruction_master_read),                       //                                                           .read
		.nios2_gen2_0_instruction_master_readdata                         (nios2_gen2_0_instruction_master_readdata),                   //                                                           .readdata
		.nios2_gen2_0_instruction_master_readdatavalid                    (nios2_gen2_0_instruction_master_readdatavalid),              //                                                           .readdatavalid
		.jtag_uart_avalon_jtag_slave_address                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //                                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                                           .write
		.jtag_uart_avalon_jtag_slave_read                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                                           .read
		.jtag_uart_avalon_jtag_slave_readdata                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                                           .chipselect
		.leds_0_s1_address                                                (mm_interconnect_0_leds_0_s1_address),                        //                                                  leds_0_s1.address
		.leds_0_s1_write                                                  (mm_interconnect_0_leds_0_s1_write),                          //                                                           .write
		.leds_0_s1_readdata                                               (mm_interconnect_0_leds_0_s1_readdata),                       //                                                           .readdata
		.leds_0_s1_writedata                                              (mm_interconnect_0_leds_0_s1_writedata),                      //                                                           .writedata
		.leds_0_s1_chipselect                                             (mm_interconnect_0_leds_0_s1_chipselect),                     //                                                           .chipselect
		.nios2_gen2_0_debug_mem_slave_address                             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //                               nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                                           .write
		.nios2_gen2_0_debug_mem_slave_read                                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                                           .read
		.nios2_gen2_0_debug_mem_slave_readdata                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                                           .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                                           .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                                           .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                                           .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                                           .debugaccess
		.onchip_memory2_0_s1_address                                      (mm_interconnect_0_onchip_memory2_0_s1_address),              //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                                           .clken
		.sdram_controller_0_s1_address                                    (mm_interconnect_0_sdram_controller_0_s1_address),            //                                      sdram_controller_0_s1.address
		.sdram_controller_0_s1_write                                      (mm_interconnect_0_sdram_controller_0_s1_write),              //                                                           .write
		.sdram_controller_0_s1_read                                       (mm_interconnect_0_sdram_controller_0_s1_read),               //                                                           .read
		.sdram_controller_0_s1_readdata                                   (mm_interconnect_0_sdram_controller_0_s1_readdata),           //                                                           .readdata
		.sdram_controller_0_s1_writedata                                  (mm_interconnect_0_sdram_controller_0_s1_writedata),          //                                                           .writedata
		.sdram_controller_0_s1_byteenable                                 (mm_interconnect_0_sdram_controller_0_s1_byteenable),         //                                                           .byteenable
		.sdram_controller_0_s1_readdatavalid                              (mm_interconnect_0_sdram_controller_0_s1_readdatavalid),      //                                                           .readdatavalid
		.sdram_controller_0_s1_waitrequest                                (mm_interconnect_0_sdram_controller_0_s1_waitrequest),        //                                                           .waitrequest
		.sdram_controller_0_s1_chipselect                                 (mm_interconnect_0_sdram_controller_0_s1_chipselect),         //                                                           .chipselect
		.sysid_control_slave_address                                      (mm_interconnect_0_sysid_control_slave_address),              //                                        sysid_control_slave.address
		.sysid_control_slave_readdata                                     (mm_interconnect_0_sysid_control_slave_readdata),             //                                                           .readdata
		.sysid_qsys_0_control_slave_address                               (mm_interconnect_0_sysid_qsys_0_control_slave_address),       //                                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)       //                                                           .readdata
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_irq_mapper_002 irq_mapper_002 (
		.clk           (pll_0_outclk0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_0_outclk0_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (pll_0_outclk1_clk),                      //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
